module x86_64

pub fn (a &Arch) initialize_early() {

}

pub fn (a &Arch) initialize() {

}