module cpu