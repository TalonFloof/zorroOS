module limine

// Implementation of the Limine Protocol Structs in V

