module panic

pub enum ZorroPanicCategory as u8 {
	generic = 1
	incompatable_hardware = 2
	out_of_memory = 3
	ramdisk = 4
}

const (
	generic_panic_img = [
		u8(0x00),0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x80,0xC0,0x00,
		0x00,0x00,0xE1,0x40,0x00,
		0x00,0x00,0x92,0x40,0x00,
		0x00,0x00,0x4E,0x40,0x00,
		0x00,0x00,0x4F,0xC0,0x00,
		0x00,0x00,0x7F,0xC0,0x00,
		0x00,0x00,0x6B,0xC0,0x00,
		0x00,0x00,0x77,0xC0,0x00,
		0x00,0x00,0xEB,0xC0,0x00,
		0x00,0x01,0xFF,0xD0,0x00,
		0x00,0x01,0xFF,0xE0,0x00,
		0x00,0x80,0x3F,0xF0,0x00,
		0x00,0xC0,0x3F,0xFC,0x00,
		0x00,0x61,0xFF,0xF8,0x00,
		0x01,0x23,0xFF,0xFC,0x00,
		0x31,0x87,0xFF,0xFE,0x00,
		0x1C,0xC7,0xFF,0xFC,0x00,
		0x06,0x27,0xBF,0xFE,0x00,
		0x00,0x83,0x1F,0xFE,0x00,
		0x00,0x0E,0x1B,0xFF,0x00,
		0x02,0xD3,0x95,0xFE,0x00,
		0x01,0x98,0xDB,0xFE,0x00,
		0x01,0x3E,0x7F,0xFF,0x00,
		0x00,0x3F,0x9F,0xFE,0x00,
		0x00,0x1F,0xDF,0xFE,0x00,
		0x00,0x0F,0xFF,0xFE,0x00,
		0x00,0x01,0xFF,0xFF,0x00,
		0x00,0x00,0xFF,0xFC,0x00,
		0x00,0x00,0xFF,0xFA,0x00,
		0x00,0x03,0xFF,0xF8,0x00,
		0x00,0x0F,0xFF,0xF8,0x00,
		0x00,0x17,0xFF,0xF0,0x00,
		0x00,0x13,0xFF,0xE0,0x00,
		0x00,0x11,0xFF,0xC0,0x00,
		0x00,0x1F,0xFF,0x80,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
	]!
	incompatable_hardware_img = [
		u8(0x00),0x04,0x00,0x00,0x00,
		0x00,0x02,0x00,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x02,0x00,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x02,0x00,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x02,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x02,0x00,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x42,0x60,0x00,0x00,
		0x00,0x70,0xA0,0x00,0x00,
		0x00,0x49,0x20,0x00,0x00,
		0x00,0x27,0x20,0x00,0x00,
		0x00,0x27,0xE0,0x00,0x00,
		0x00,0x3F,0xE4,0x00,0x00,
		0x00,0x39,0xF8,0x00,0x00,
		0x00,0x35,0xF0,0x00,0x00,
		0x00,0x73,0xFA,0x00,0x00,
		0x00,0xFF,0xFC,0x00,0x00,
		0xC0,0xFF,0xFA,0x00,0x00,
		0xF0,0x0F,0xFC,0x80,0x00,
		0xFC,0x0F,0xFF,0x00,0x00,
		0xFF,0x0F,0xFE,0x00,0x00,
		0xFF,0xCF,0xFF,0x40,0x00,
		0xFF,0xEF,0xFF,0x80,0x00,
		0xFF,0xEF,0xFF,0x10,0x00,
		0xFF,0x2F,0xFF,0xA0,0x00,
		0xFC,0x2F,0xFF,0xC0,0x00,
		0xF1,0xAF,0xFF,0xE8,0x00,
		0xC6,0xAF,0xFF,0xF0,0x00,
		0x98,0xA7,0xFF,0xE0,0xE0,
		0xAA,0xA7,0xFF,0xE9,0x20,
		0xA0,0xA7,0xFF,0xF2,0x20,
		0xA4,0xA7,0xFF,0xF7,0x40,
		0xAA,0xA7,0xFF,0xF7,0x80,
		0xA0,0xA7,0xFF,0xFF,0x00,
		0xA1,0xA7,0xFF,0xFF,0x00,
		0xA6,0x27,0xFF,0xFE,0x00,
		0xB8,0x27,0xFF,0xFC,0x00,
		0x80,0x27,0xFF,0xE0,0x00,
		0x80,0x23,0xFF,0xC0,0x00,
		0x80,0x20,0x00,0x00,0x00,
		0x80,0xC0,0x00,0x00,0x00,
	]!
	out_of_memory_img = [
		u8(0x00),0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x04,0x00,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x09,0x00,0x00,0x00,
		0x00,0x0A,0x00,0x00,0x00,
		0x00,0x42,0x60,0x00,0x00,
		0x00,0x70,0xA0,0x00,0x00,
		0x00,0x49,0x20,0x00,0x00,
		0x00,0x27,0x20,0x00,0x00,
		0x00,0x27,0xE0,0x00,0x00,
		0x00,0x3F,0xE0,0x00,0x00,
		0x00,0x3D,0xF0,0x00,0x00,
		0x00,0x39,0xF0,0x00,0x00,
		0x00,0x73,0xF8,0x00,0x00,
		0x00,0xFF,0xF8,0x00,0x00,
		0x00,0xFF,0xF8,0x00,0x00,
		0x00,0x0F,0xFC,0x00,0x00,
		0x00,0x0F,0xFE,0x00,0x00,
		0x00,0x0F,0xFE,0x00,0x00,
		0x00,0x0F,0xFF,0x00,0x00,
		0x00,0x0F,0xFF,0x00,0x00,
		0x00,0xFF,0xFF,0x00,0x00,
		0x01,0xFF,0xFF,0x80,0x00,
		0x0D,0xFF,0xFF,0xC0,0x00,
		0x33,0xCF,0xFF,0xE0,0x00,
		0x40,0x8F,0xFF,0xE0,0x00,
		0x73,0x87,0xFF,0xE0,0xE0,
		0xCC,0xC7,0xFF,0xE1,0x20,
		0x40,0xA7,0xFF,0xF2,0x20,
		0xB3,0x67,0xFF,0xF7,0x40,
		0x4C,0x67,0xFF,0xF7,0x80,
		0xA2,0xA7,0xFF,0xFF,0x00,
		0x55,0x67,0xFF,0xFF,0x00,
		0xAA,0xA7,0xFF,0xFE,0x00,
		0x55,0x67,0xFF,0xFC,0x00,
		0xAA,0xA7,0xFF,0xE0,0x00,
		0x55,0x63,0xFF,0xC0,0x00,
		0xAA,0xA0,0x00,0x00,0x00,
		0x55,0x60,0x00,0x00,0x00,
	]!
	ramdisk_img = [
		u8(0x00),0x0A,0x00,0x00,0x00,
		0x00,0x15,0x00,0x00,0x00,
		0x00,0x0A,0x80,0x00,0x00,
		0x00,0x11,0x00,0x00,0x00,
		0x00,0x00,0x80,0x00,0x00,
		0x00,0x01,0x00,0x00,0x00,
		0x00,0x02,0x80,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x00,0x00,0x00,0x00,
		0x00,0x02,0x00,0x00,0x00,
		0x00,0x05,0x00,0x00,0x00,
		0x00,0x42,0x60,0x00,0x00,
		0x00,0x70,0xA0,0x00,0x00,
		0x00,0x49,0x20,0x00,0x00,
		0x00,0x27,0x20,0x00,0x00,
		0x00,0x27,0xE0,0x00,0x00,
		0x00,0x3F,0xE0,0x00,0x00,
		0x00,0x3D,0xF0,0x00,0x00,
		0x00,0x33,0xF0,0x00,0x00,
		0x00,0x7F,0xF8,0x00,0x00,
		0x00,0xFF,0xF8,0x00,0x00,
		0x00,0xFF,0xF8,0x00,0x00,
		0x00,0x0F,0xFC,0x00,0x00,
		0x00,0x0F,0xFE,0x00,0x00,
		0x00,0x0F,0xFE,0x00,0x00,
		0x00,0x0F,0xFF,0x00,0x00,
		0x00,0x0F,0xFF,0x00,0x00,
		0x60,0x0F,0xFF,0x00,0x00,
		0xF8,0x0F,0xFF,0x80,0x00,
		0xFE,0x0F,0xFF,0xC0,0x00,
		0xFF,0x8F,0xFF,0xE0,0x00,
		0xF9,0xEF,0xFF,0xE0,0x00,
		0xE6,0x77,0xFF,0xE0,0xE0,
		0xDF,0xB7,0xFF,0xE1,0x20,
		0xDF,0xB7,0xFF,0xF2,0x20,
		0xB9,0xD7,0xFF,0xF7,0x40,
		0xB9,0xD7,0xFF,0xF7,0x80,
		0xDF,0xB7,0xFF,0xFF,0x00,
		0xDF,0xA7,0xFF,0xFF,0x00,
		0xE6,0x47,0xFF,0xFE,0x00,
		0x79,0x97,0xFF,0xFC,0x00,
		0x1F,0x37,0xFF,0xE0,0x00,
		0x06,0x73,0xFF,0xC0,0x00,
		0x00,0xF0,0x00,0x00,0x00,
		0x00,0x60,0x00,0x00,0x00,
	]!
)

[noreturn]
pub fn panic_multiline(category ZorroPanicCategory, msg &string, len int) {
	log := zorro_arch.get_logger() or { unsafe { goto panic_framebuffer } return}
	if category != .ramdisk {
		log.fatal("Kernel Panic (hart 0x0)")
		log.fatal(msg)
	}
panic_framebuffer:
	fb := zorro_arch.get_framebuffer() or { unsafe { goto panic_halt } return }
	res := fb.get_resolution()
	for y in 0 .. res.h { // Dim Screen
		for x in 0 .. res.w {
			fb.set(x,y,(fb.get(x,y) >> 1) & 0x7f7f7f7f)
		}
	}
	match category {
		.generic {
			fb.render_monochrome_bitmap(int(res.w)/2-(35*3/2),int(res.h)/2-(45*3/2),35,45,3,0xffffff,5,&generic_panic_img)
		}
		.incompatable_hardware {
			fb.render_monochrome_bitmap(int(res.w)/2-(35*3/2),int(res.h)/2-(45*3/2),35,45,3,0xffffff,5,&incompatable_hardware_img)
		}
		.out_of_memory {
			fb.render_monochrome_bitmap(int(res.w)/2-(35*3/2),int(res.h)/2-(45*3/2),35,45,3,0xffffff,5,&out_of_memory_img)
		}
		.ramdisk {
			fb.render_monochrome_bitmap(int(res.w)/2-(35*3/2),int(res.h)/2-(45*3/2),35,45,3,0xffffff,5,&ramdisk_img)
		}
	}
	if category != .ramdisk {
		fb.draw_centered_text_literal(int(res.w)/2,int(res.h)/2+(45*3/2),1,0xffffff,"Kernel Panic")
		for i := 0; i < len; i++ {
			unsafe {
				fb.draw_centered_text(int(res.w)/2,(int(res.h)/2+(45*3/2))+16+(i*16),1,0xffffff,&(msg[i]))
			}
		}
	} else {
		for i := 0; i < len; i++ {
			unsafe {
				fb.draw_centered_text(int(res.w)/2,int(res.h)/2+(45*3/2)+(i*16),1,0xffffff,&(msg[i]))
			}
		}
	}
panic_halt:
	zorro_arch.halt()
}

[export: "kpanic"]
[noreturn]
pub fn panic(category ZorroPanicCategory, msg string) {
	panic_multiline(category,&msg,1)
}