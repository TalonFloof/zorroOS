module framebuffer_impl

