module framebuffer

pub struct ZorroFramebufferResolution {
pub:
	w int
	h int
}

pub interface IZorroFramebuffer {
	get_resolution() ZorroFramebufferResolution
	get_depth() u8
	get(int,int) u32
	get_unsafe_pointer() &u8
	set(int,int,u32)
}

pub fn (fb &IZorroFramebuffer) rect(x int, y int, w int, h int, color u32) {
	for i in y .. (y+h) {
		for j in x .. (x+w) {
			fb.set(j,i,color)
		}
	}
}

pub fn (fb &IZorroFramebuffer) clear(color u32) {
	resolution := fb.get_resolution()
	fb.rect(0,0,resolution.w,resolution.h,color)
}

pub fn (fb &IZorroFramebuffer) render_monochrome_bitmap(x int, y int, w int, h int, scale int, color u32, line_size u64, ptr &u8) {
	for i in 0 .. h {
		for j in 0 .. w {
			byte_offset := (u64(i)*line_size)+(u64(j)/8)
			bit_offset := u64(j) % 8
			dat := unsafe {ptr[byte_offset]}
			if dat & (1 << (7-bit_offset)) != 0 {
				fb.rect(x+(j*scale),y+(i*scale),scale,scale,color)
			}
		}
	}
}

const (
	zorro_script = [u8(170), 0, 128, 0, 128, 74, 234, 90, 201, 0, 128, 0, 128, 0, 128, 85, 170,
		0, 128, 0, 128, 57, 194, 50, 138, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 59,
		193, 49, 137, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 123, 193, 121, 193, 121,
		128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 121, 194, 122, 194, 121, 128, 0, 128, 0,
		128, 85, 170, 0, 128, 0, 128, 122, 194, 123, 194, 122, 128, 0, 128, 0, 128, 85, 170, 0,
		128, 0, 128, 49, 202, 122, 202, 73, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 115,
		202, 115, 202, 115, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 30, 145, 30, 145, 30,
		128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 34, 162, 62, 162, 34, 128, 0, 128, 0, 128,
		85, 170, 0, 128, 0, 128, 32, 160, 32, 160, 62, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0,
		128, 34, 162, 34, 148, 8, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 62, 160, 62, 160,
		32, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 30, 160, 32, 160, 30, 128, 0, 128, 0,
		128, 85, 170, 0, 128, 0, 128, 30, 160, 28, 130, 60, 128, 0, 128, 0, 128, 85, 170, 0, 128,
		0, 128, 30, 160, 28, 130, 60, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 57, 165, 37,
		165, 57, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 113, 202, 74, 202, 113, 128, 0,
		128, 0, 128, 85, 170, 0, 128, 0, 128, 113, 202, 74, 202, 113, 128, 0, 128, 0, 128, 85,
		170, 0, 128, 0, 128, 113, 202, 74, 202, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128,
		113, 202, 74, 202, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 73, 234, 106, 219,
		74, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 52, 194, 49, 137, 113, 128, 0, 128, 0,
		128, 85, 170, 0, 128, 0, 128, 123, 193, 121, 193, 121, 128, 0, 128, 0, 128, 85, 170, 0,
		128, 0, 128, 51, 196, 71, 196, 52, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 62, 160,
		62, 160, 62, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 58, 194, 50, 138, 113, 128,
		0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 121, 194, 121, 192, 123, 128, 0, 128, 0, 128,
		85, 170, 0, 128, 0, 128, 30, 144, 30, 144, 16, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0,
		128, 14, 144, 22, 146, 14, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 28, 146, 28, 148,
		18, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 18, 146, 18, 146, 12, 128, 0, 128, 0,
		128, 85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 8, 8, 8, 8,
		8, 0, 8, 8, 0, 0, 0, 0, 34, 34, 34, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 18,
		18, 126, 36, 36, 126, 72, 72, 72, 0, 0, 0, 0, 0, 0, 8, 62, 73, 72, 56, 14, 9, 73, 62, 8,
		0, 0, 0, 0, 0, 0, 49, 74, 74, 52, 8, 8, 22, 41, 41, 70, 0, 0, 0, 0, 0, 0, 28, 34, 34, 20,
		24, 41, 69, 66, 70, 57, 0, 0, 0, 0, 8, 8, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		4, 8, 8, 16, 16, 16, 16, 16, 16, 8, 8, 4, 0, 0, 0, 0, 32, 16, 16, 8, 8, 8, 8, 8, 8, 16,
		16, 32, 0, 0, 0, 0, 0, 0, 0, 8, 73, 42, 28, 42, 73, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8,
		8, 127, 8, 8, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 8, 8, 16, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 24, 0, 0,
		0, 0, 0, 0, 2, 2, 4, 8, 8, 16, 16, 32, 64, 64, 0, 0, 0, 0, 0, 0, 24, 36, 66, 70, 74, 82,
		98, 66, 36, 24, 0, 0, 0, 0, 0, 0, 8, 24, 40, 8, 8, 8, 8, 8, 8, 62, 0, 0, 0, 0, 0, 0, 60,
		66, 66, 2, 12, 16, 32, 64, 64, 126, 0, 0, 0, 0, 0, 0, 60, 66, 66, 2, 28, 2, 2, 66, 66,
		60, 0, 0, 0, 0, 0, 0, 4, 12, 20, 36, 68, 68, 126, 4, 4, 4, 0, 0, 0, 0, 0, 0, 126, 64, 64,
		64, 124, 2, 2, 2, 66, 60, 0, 0, 0, 0, 0, 0, 28, 32, 64, 64, 124, 66, 66, 66, 66, 60, 0,
		0, 0, 0, 0, 0, 126, 2, 2, 4, 4, 4, 8, 8, 8, 8, 0, 0, 0, 0, 0, 0, 60, 66, 66, 66, 60, 66,
		66, 66, 66, 60, 0, 0, 0, 0, 0, 0, 60, 66, 66, 66, 62, 2, 2, 2, 4, 56, 0, 0, 0, 0, 0, 0,
		0, 0, 24, 24, 0, 0, 0, 24, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 24, 0, 0, 0, 24, 8, 8, 16,
		0, 0, 0, 0, 0, 0, 2, 4, 8, 16, 32, 16, 8, 4, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 126, 0, 0, 0,
		126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 32, 16, 8, 4, 8, 16, 32, 64, 0, 0, 0, 0, 0, 0, 60,
		66, 66, 2, 4, 8, 8, 0, 8, 8, 0, 0, 0, 0, 0, 0, 28, 34, 74, 86, 82, 82, 82, 78, 32, 30,
		0, 0, 0, 0, 0, 0, 24, 36, 36, 66, 66, 126, 66, 66, 66, 66, 0, 0, 0, 0, 0, 0, 124, 66, 66,
		66, 124, 66, 66, 66, 66, 124, 0, 0, 0, 0, 0, 0, 60, 66, 66, 64, 64, 64, 64, 66, 66, 60,
		0, 0, 0, 0, 0, 0, 120, 68, 66, 66, 66, 66, 66, 66, 68, 120, 0, 0, 0, 0, 0, 0, 126, 64,
		64, 64, 124, 64, 64, 64, 64, 126, 0, 0, 0, 0, 0, 0, 126, 64, 64, 64, 124, 64, 64, 64, 64,
		64, 0, 0, 0, 0, 0, 0, 60, 66, 66, 64, 64, 78, 66, 66, 70, 58, 0, 0, 0, 0, 0, 0, 66, 66,
		66, 66, 126, 66, 66, 66, 66, 66, 0, 0, 0, 0, 0, 0, 62, 8, 8, 8, 8, 8, 8, 8, 8, 62, 0, 0,
		0, 0, 0, 0, 31, 4, 4, 4, 4, 4, 4, 68, 68, 56, 0, 0, 0, 0, 0, 0, 66, 68, 72, 80, 96, 96,
		80, 72, 68, 66, 0, 0, 0, 0, 0, 0, 64, 64, 64, 64, 64, 64, 64, 64, 64, 126, 0, 0, 0, 0,
		0, 0, 66, 66, 102, 102, 90, 90, 66, 66, 66, 66, 0, 0, 0, 0, 0, 0, 66, 98, 98, 82, 82, 74,
		74, 70, 70, 66, 0, 0, 0, 0, 0, 0, 60, 66, 66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 0, 0, 0,
		0, 124, 66, 66, 66, 124, 64, 64, 64, 64, 64, 0, 0, 0, 0, 0, 0, 60, 66, 66, 66, 66, 66,
		66, 90, 102, 60, 3, 0, 0, 0, 0, 0, 124, 66, 66, 66, 124, 72, 68, 68, 66, 66, 0, 0, 0, 0,
		0, 0, 60, 66, 66, 64, 48, 12, 2, 66, 66, 60, 0, 0, 0, 0, 0, 0, 127, 8, 8, 8, 8, 8, 8, 8,
		8, 8, 0, 0, 0, 0, 0, 0, 66, 66, 66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 0, 0, 0, 0, 65, 65,
		65, 34, 34, 34, 20, 20, 8, 8, 0, 0, 0, 0, 0, 0, 66, 66, 66, 66, 90, 90, 102, 102, 66, 66,
		0, 0, 0, 0, 0, 0, 66, 66, 36, 36, 24, 24, 36, 36, 66, 66, 0, 0, 0, 0, 0, 0, 65, 65, 34,
		34, 20, 8, 8, 8, 8, 8, 0, 0, 0, 0, 0, 0, 126, 2, 2, 4, 8, 16, 32, 64, 64, 126, 0, 0, 0,
		0, 0, 14, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 14, 0, 0, 0, 0, 0, 64, 64, 32, 16, 16, 8, 8, 4,
		2, 2, 0, 0, 0, 0, 0, 112, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 112, 0, 0, 0, 24, 36,
		66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 127, 0,
		0, 32, 16, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 66, 2, 62, 66,
		66, 70, 58, 0, 0, 0, 0, 0, 64, 64, 64, 92, 98, 66, 66, 66, 66, 98, 92, 0, 0, 0, 0, 0, 0,
		0, 0, 60, 66, 64, 64, 64, 64, 66, 60, 0, 0, 0, 0, 0, 2, 2, 2, 58, 70, 66, 66, 66, 66, 70,
		58, 0, 0, 0, 0, 0, 0, 0, 0, 60, 66, 66, 126, 64, 64, 66, 60, 0, 0, 0, 0, 0, 12, 16, 16,
		16, 124, 16, 16, 16, 16, 16, 16, 0, 0, 0, 0, 0, 0, 0, 2, 58, 68, 68, 68, 56, 32, 60, 66,
		66, 60, 0, 0, 0, 64, 64, 64, 92, 98, 66, 66, 66, 66, 66, 66, 0, 0, 0, 0, 0, 8, 8, 0, 24,
		8, 8, 8, 8, 8, 8, 62, 0, 0, 0, 0, 0, 4, 4, 0, 12, 4, 4, 4, 4, 4, 4, 4, 72, 48, 0, 0, 0,
		64, 64, 64, 68, 72, 80, 96, 80, 72, 68, 66, 0, 0, 0, 0, 0, 24, 8, 8, 8, 8, 8, 8, 8, 8,
		8, 62, 0, 0, 0, 0, 0, 0, 0, 0, 118, 73, 73, 73, 73, 73, 73, 73, 0, 0, 0, 0, 0, 0, 0, 0,
		92, 98, 66, 66, 66, 66, 66, 66, 0, 0, 0, 0, 0, 0, 0, 0, 60, 66, 66, 66, 66, 66, 66, 60,
		0, 0, 0, 0, 0, 0, 0, 0, 92, 98, 66, 66, 66, 66, 98, 92, 64, 64, 0, 0, 0, 0, 0, 0, 58, 70,
		66, 66, 66, 66, 70, 58, 2, 2, 0, 0, 0, 0, 0, 0, 92, 98, 66, 64, 64, 64, 64, 64, 0, 0, 0,
		0, 0, 0, 0, 0, 60, 66, 64, 48, 12, 2, 66, 60, 0, 0, 0, 0, 0, 0, 16, 16, 16, 124, 16, 16,
		16, 16, 16, 12, 0, 0, 0, 0, 0, 0, 0, 0, 66, 66, 66, 66, 66, 66, 70, 58, 0, 0, 0, 0, 0,
		0, 0, 0, 66, 66, 66, 36, 36, 36, 24, 24, 0, 0, 0, 0, 0, 0, 0, 0, 65, 73, 73, 73, 73, 73,
		73, 54, 0, 0, 0, 0, 0, 0, 0, 0, 66, 66, 36, 24, 24, 36, 66, 66, 0, 0, 0, 0, 0, 0, 0, 0,
		66, 66, 66, 66, 66, 38, 26, 2, 2, 60, 0, 0, 0, 0, 0, 0, 126, 2, 4, 8, 16, 32, 64, 126,
		0, 0, 0, 0, 0, 12, 16, 16, 8, 8, 16, 32, 16, 8, 8, 16, 16, 12, 0, 0, 8, 8, 8, 8, 8, 8,
		8, 8, 8, 8, 8, 8, 8, 8, 0, 0, 0, 48, 8, 8, 16, 16, 8, 4, 8, 16, 16, 8, 8, 48, 0, 0, 0,
		49, 73, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 128, 0, 128, 115, 202, 75, 202, 115,
		128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 113, 202, 115, 194, 66, 128, 0, 128, 0, 128,
		85, 170, 0, 128, 0, 128, 73, 202, 122, 202, 73, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0,
		128, 115, 202, 115, 202, 114, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 75, 234, 91,
		202, 75, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 116, 166, 37, 164, 116, 128, 0,
		128, 0, 128, 85, 170, 0, 128, 0, 128, 75, 234, 91, 202, 75, 128, 0, 128, 0, 128, 85, 170,
		0, 128, 0, 128, 57, 194, 49, 136, 115, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 121,
		194, 121, 192, 123, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 75, 201, 121, 201, 73,
		128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 37, 164, 60, 164, 36, 128, 0, 128, 0, 128,
		85, 170, 0, 128, 0, 128, 69, 196, 68, 168, 16, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0,
		128, 114, 202, 114, 194, 67, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 114, 202, 114,
		194, 67, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 14, 137, 14, 138, 9, 128, 0, 128,
		0, 128, 85, 170, 0, 128, 0, 128, 57, 194, 49, 136, 115, 128, 0, 128, 0, 128, 85, 170, 0,
		128, 0, 128, 57, 194, 49, 136, 115, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 113,
		202, 74, 202, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 114, 202, 114, 194, 65,
		128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 114, 202, 114, 194, 65, 128, 0, 128, 0, 128,
		85, 170, 0, 128, 0, 128, 59, 193, 49, 137, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0,
		128, 57, 194, 66, 194, 57, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 34, 182, 42, 162,
		34, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 59, 194, 51, 138, 114, 128, 0, 128, 0,
		128, 85, 170, 0, 128, 0, 128, 123, 194, 123, 194, 122, 128, 0, 128, 0, 128, 85, 170, 0,
		128, 0, 128, 57, 194, 50, 138, 113, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 51, 196,
		37, 148, 99, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 57, 194, 50, 138, 113, 128,
		0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 57, 194, 65, 192, 59, 128, 0, 128, 0, 128, 85,
		170, 0, 128, 0, 128, 14, 144, 12, 130, 28, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128,
		49, 202, 73, 200, 51, 128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 28, 146, 28, 144, 16,
		128, 0, 128, 0, 128, 85, 170, 0, 128, 0, 128, 51, 202, 123, 202, 74, 128, 0, 128, 0, 128,
		85, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 8, 8, 8, 8, 8,
		8, 8, 0, 0, 0, 0, 0, 0, 8, 8, 62, 73, 72, 72, 73, 62, 8, 8, 0, 0, 0, 0, 0, 0, 14, 16, 16,
		16, 124, 16, 16, 16, 62, 97, 0, 0, 0, 0, 0, 0, 0, 66, 60, 36, 66, 66, 36, 60, 66, 0, 0,
		0, 0, 0, 0, 0, 65, 34, 20, 8, 127, 8, 127, 8, 8, 8, 0, 0, 0, 0, 0, 0, 8, 8, 8, 8, 0, 0,
		8, 8, 8, 8, 0, 0, 0, 0, 0, 0, 60, 66, 64, 60, 66, 66, 60, 2, 66, 60, 0, 0, 36, 36, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 66, 153, 165, 161, 161, 165, 153, 66,
		60, 0, 0, 0, 0, 28, 2, 30, 34, 30, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 18, 36,
		36, 72, 36, 36, 18, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 126, 2, 2, 2, 0, 0, 170, 0,
		128, 58, 194, 51, 138, 114, 128, 0, 128, 3, 128, 0, 128, 85, 0, 0, 0, 0, 60, 66, 185, 165,
		165, 185, 169, 165, 66, 60, 0, 0, 0, 0, 126, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 24, 36, 36, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 8, 127, 8, 8, 8, 0,
		127, 0, 0, 0, 0, 0, 0, 56, 68, 4, 24, 32, 64, 124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 68, 4,
		56, 4, 68, 56, 0, 0, 0, 0, 0, 0, 0, 4, 8, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 66, 66, 66, 66, 66, 66, 102, 89, 64, 128, 0, 0, 0, 0, 63, 122, 122, 122, 58,
		10, 10, 10, 10, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 48, 0, 0, 0, 16, 48, 80, 16, 16, 16, 124, 0, 0, 0, 0,
		0, 0, 0, 0, 28, 34, 34, 34, 28, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 72, 36,
		36, 18, 36, 36, 72, 72, 0, 0, 0, 0, 0, 0, 34, 98, 36, 40, 40, 18, 22, 42, 78, 66, 0, 0,
		0, 0, 0, 0, 34, 98, 36, 40, 40, 20, 26, 34, 68, 78, 0, 0, 0, 0, 0, 0, 98, 18, 36, 24, 104,
		18, 22, 42, 78, 66, 0, 0, 0, 0, 0, 0, 16, 16, 0, 16, 16, 32, 64, 66, 66, 60, 0, 0, 48,
		12, 0, 0, 24, 36, 36, 66, 66, 126, 66, 66, 66, 66, 0, 0, 12, 48, 0, 0, 24, 36, 36, 66,
		66, 126, 66, 66, 66, 66, 0, 0, 24, 36, 0, 0, 24, 36, 36, 66, 66, 126, 66, 66, 66, 66, 0,
		0, 50, 76, 0, 0, 24, 36, 36, 66, 66, 126, 66, 66, 66, 66, 0, 0, 36, 36, 0, 0, 24, 36, 36,
		66, 66, 126, 66, 66, 66, 66, 0, 0, 24, 36, 24, 0, 24, 36, 36, 66, 66, 126, 66, 66, 66,
		66, 0, 0, 0, 0, 0, 0, 31, 40, 72, 72, 127, 72, 72, 72, 72, 79, 0, 0, 0, 0, 0, 0, 60, 66,
		66, 64, 64, 64, 64, 66, 66, 60, 8, 48, 48, 12, 0, 0, 126, 64, 64, 64, 124, 64, 64, 64,
		64, 126, 0, 0, 12, 48, 0, 0, 126, 64, 64, 64, 124, 64, 64, 64, 64, 126, 0, 0, 24, 36, 0,
		0, 126, 64, 64, 64, 124, 64, 64, 64, 64, 126, 0, 0, 36, 36, 0, 0, 126, 64, 64, 64, 124,
		64, 64, 64, 64, 126, 0, 0, 24, 6, 0, 0, 62, 8, 8, 8, 8, 8, 8, 8, 8, 62, 0, 0, 12, 48, 0,
		0, 62, 8, 8, 8, 8, 8, 8, 8, 8, 62, 0, 0, 24, 36, 0, 0, 62, 8, 8, 8, 8, 8, 8, 8, 8, 62,
		0, 0, 36, 36, 0, 0, 62, 8, 8, 8, 8, 8, 8, 8, 8, 62, 0, 0, 0, 0, 0, 0, 120, 68, 66, 66,
		242, 66, 66, 66, 68, 120, 0, 0, 50, 76, 0, 0, 66, 98, 98, 82, 82, 74, 74, 70, 70, 66, 0,
		0, 48, 12, 0, 0, 60, 66, 66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 12, 48, 0, 0, 60, 66, 66,
		66, 66, 66, 66, 66, 66, 60, 0, 0, 24, 36, 0, 0, 60, 66, 66, 66, 66, 66, 66, 66, 66, 60,
		0, 0, 50, 76, 0, 0, 60, 66, 66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 36, 36, 0, 0, 60, 66,
		66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66, 36, 24, 36, 66, 0, 0, 0,
		0, 0, 0, 0, 2, 58, 68, 70, 74, 74, 82, 82, 98, 34, 92, 64, 0, 48, 12, 0, 0, 66, 66, 66,
		66, 66, 66, 66, 66, 66, 60, 0, 0, 12, 48, 0, 0, 66, 66, 66, 66, 66, 66, 66, 66, 66, 60,
		0, 0, 24, 36, 0, 0, 66, 66, 66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 36, 36, 0, 0, 66, 66,
		66, 66, 66, 66, 66, 66, 66, 60, 0, 0, 12, 48, 0, 0, 65, 65, 34, 34, 20, 8, 8, 8, 8, 8,
		0, 0, 0, 0, 0, 64, 64, 120, 68, 66, 66, 68, 120, 64, 64, 64, 0, 0, 0, 0, 0, 0, 56, 68,
		68, 72, 88, 68, 66, 66, 82, 76, 0, 0, 0, 0, 48, 12, 0, 0, 60, 66, 2, 62, 66, 66, 70, 58,
		0, 0, 0, 0, 12, 48, 0, 0, 60, 66, 2, 62, 66, 66, 70, 58, 0, 0, 0, 0, 24, 36, 0, 0, 60,
		66, 2, 62, 66, 66, 70, 58, 0, 0, 0, 0, 50, 76, 0, 0, 60, 66, 2, 62, 66, 66, 70, 58, 0,
		0, 0, 0, 36, 36, 0, 0, 60, 66, 2, 62, 66, 66, 70, 58, 0, 0, 0, 24, 36, 24, 0, 0, 60, 66,
		2, 62, 66, 66, 70, 58, 0, 0, 0, 0, 0, 0, 0, 0, 62, 73, 9, 63, 72, 72, 73, 62, 0, 0, 0,
		0, 0, 0, 0, 0, 60, 66, 64, 64, 64, 64, 66, 60, 8, 48, 0, 0, 48, 12, 0, 0, 60, 66, 66, 126,
		64, 64, 66, 60, 0, 0, 0, 0, 12, 48, 0, 0, 60, 66, 66, 126, 64, 64, 66, 60, 0, 0, 0, 0,
		24, 36, 0, 0, 60, 66, 66, 126, 64, 64, 66, 60, 0, 0, 0, 0, 36, 36, 0, 0, 60, 66, 66, 126,
		64, 64, 66, 60, 0, 0, 0, 0, 48, 12, 0, 0, 24, 8, 8, 8, 8, 8, 8, 62, 0, 0, 0, 0, 12, 48,
		0, 0, 24, 8, 8, 8, 8, 8, 8, 62, 0, 0, 0, 0, 24, 36, 0, 0, 24, 8, 8, 8, 8, 8, 8, 62, 0,
		0, 0, 0, 36, 36, 0, 0, 24, 8, 8, 8, 8, 8, 8, 62, 0, 0, 0, 0, 50, 12, 20, 34, 2, 62, 66,
		66, 66, 66, 66, 60, 0, 0, 0, 0, 50, 76, 0, 0, 92, 98, 66, 66, 66, 66, 66, 66, 0, 0, 0,
		0, 48, 12, 0, 0, 60, 66, 66, 66, 66, 66, 66, 60, 0, 0, 0, 0, 12, 48, 0, 0, 60, 66, 66,
		66, 66, 66, 66, 60, 0, 0, 0, 0, 24, 36, 0, 0, 60, 66, 66, 66, 66, 66, 66, 60, 0, 0, 0,
		0, 50, 76, 0, 0, 60, 66, 66, 66, 66, 66, 66, 60, 0, 0, 0, 0, 36, 36, 0, 0, 60, 66, 66,
		66, 66, 66, 66, 60, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 0, 126, 0, 0, 24, 0, 0, 0, 0, 0, 0,
		0, 0, 2, 60, 70, 74, 74, 82, 82, 98, 60, 64, 0, 0, 0, 48, 12, 0, 0, 66, 66, 66, 66, 66,
		66, 70, 58, 0, 0, 0, 0, 12, 48, 0, 0, 66, 66, 66, 66, 66, 66, 70, 58, 0, 0, 0, 0, 24, 36,
		0, 0, 66, 66, 66, 66, 66, 66, 70, 58, 0, 0, 0, 0, 36, 36, 0, 0, 66, 66, 66, 66, 66, 66,
		70, 58, 0, 0, 0, 0, 12, 48, 0, 0, 66, 66, 66, 66, 66, 38, 26, 2, 2, 60, 0, 0, 0, 64, 64,
		64, 92, 98, 66, 66, 66, 66, 98, 92, 64, 64, 0, 0, 36, 36, 0, 0, 66, 66, 66, 66, 66, 38,
		26, 2, 2, 60]!
)

pub fn (fb &IZorroFramebuffer) render_rune(x int, y int, scale int, color u32, rune_ rune) {
	if u32(rune_) > 255 {
		panic("Attempted to render a rune outside of the ZorroScript font range")
	}
	fb.render_monochrome_bitmap(x,y,8,16,scale,color,1,&u8(u64(&zorro_script)+(u64(rune_)*16)))
}

pub fn (fb &IZorroFramebuffer) draw_text(x int, y int, scale int, color u32, str &string) {
	for i := 0; i < str.len; i++ {
		fb.render_rune(x+(i*(8*scale)),y,scale,color,unsafe {rune(str.str[i])})
	}
}

pub fn (fb &IZorroFramebuffer) draw_text_literal(x int, y int, scale int, color u32, str string) {
	fb.draw_text(x,y,scale,color,&str)
}

pub fn (fb &IZorroFramebuffer) draw_centered_text(center_x int, y int, scale int, color u32, str &string) {
	fb.draw_text(center_x-((str.len*(8*scale))/2),y,scale,color,str)
}

pub fn (fb &IZorroFramebuffer) draw_centered_text_literal(center_x int, y int, scale int, color u32, str string) {
	fb.draw_text(center_x-((str.len*(8*scale))/2),y,scale,color,&str)
}