module paging

pub interface VMSpace {
	
}