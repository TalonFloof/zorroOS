module logger

import arch.interfaces.logger as i_log

