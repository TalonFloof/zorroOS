module x86_64

import limine

pub fn zorro_arch_initialize() {

}