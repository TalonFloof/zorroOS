module ksync

pub struct Atomic<T> {
	
}

