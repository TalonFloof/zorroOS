module paging

