module alloc

