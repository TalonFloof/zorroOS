module paging

module paging

pub interface VMSpace {
	
}